module instructionMemory (
  input logic [31:0] Address,  
  //input logic WriteEnable,
  output logic [31:0] InstructionOut
);

logic [3:0][7:0] RegisterA [31:0];

initial begin

  RegisterA[0] = 32'b0000000_00000_00010_000_11111_0110011; // reg0,reg4,reg31,add
  RegisterA[1] = 32'b0100000_00111_00011_000_11110_0110011; // reg7,reg3,reg30,sub
  RegisterA[2] = 32'b0000000_00111_00000_001_11101_0110011; // reg7,reg0,reg29, SLL
  RegisterA[3] = 32'b0000000_00000_00100_010_11100_0110011; // reg0,reg,reg28, SLT
  RegisterA[4] = 32'b0000000_00001_00000_011_11011_0110011; // reg1,reg,reg27,SLTU
  RegisterA[5] = 32'b0000000_10100_11001_100_11010_0110011; // reg20,reg25,reg26 ,XOR
  RegisterA[6] = 32'b0000000_00011_00000_101_11001_0110011; // reg3,reg0,reg25, SRL
  RegisterA[7] = 32'b0100000_00111_00000_101_11000_0110011; // reg7,reg0,reg24, SRA
  RegisterA[8] = 32'b0000000_10100_10000_110_10111_0110011; // reg20,reg16,reg23, OR
  RegisterA[9] = 32'b0000000_10100_00001_111_10110_0110011; // reg20,reg1,reg22,AND
  
  
  RegisterA[10] = 32'b000000000101_00001_000_10110_0010011; // ,addi
  RegisterA[11] = 32'b000000000001_00010_000_10101_0010011; // ,addi
  RegisterA[12] = 32'b000000000001_00100_010_10100_0010011; // ,SLTi
  RegisterA[13] = 32'b000000000001_00100_011_10011_0010011; // ,SLTiu
  RegisterA[14] = 32'b000000000001_00100_100_10010_0010011; // ,XORi
  RegisterA[15] = 32'b000000000001_00100_110_10001_0010011; // ,ORi
  RegisterA[16] = 32'b000000000011_00010_111_10000_0010011; // ,ANDi
  RegisterA[17] = 32'b0000000_00011_00010_001_01111_0010011; // ,SLLi
  RegisterA[18] = 32'b0000000_00011_00010_101_01110_0010011; // ,SRLi
  RegisterA[19] = 32'b0000000_00011_00010_101_01101_0010011; // ,SRAi
  
    
  RegisterA[20] = 32'b000000000101_00001_000_11111_0010011; // ,addi  
  
  
  RegisterA[21] = 32'b000000000000_00001_000_01100_0000011; // ,LB
  RegisterA[22] = 32'b000000000001_00001_001_01011_0000011; // ,LH
  RegisterA[23] = 32'b000000000000_00001_010_01010_0000011; // ,LW
  RegisterA[24] = 32'b000000000000_00001_100_01001_0000011; // ,LBU
  RegisterA[25] = 32'b000000000000_00001_101_01000_0000011; // ,LHU
  
  
  RegisterA[26] = 32'b0000000_00010_00100_000_00001_0100011; //SB
  RegisterA[27] = 32'b0000000_00010_00101_001_00010_0100011; //SH
  RegisterA[28] = 32'b0000000_00010_00110_010_00011_0100011; //SW
  
  /**
  RegisterA[26] = 32'b0000000_00111_00100_000_00111_0110011; // j EXIT
  RegisterA[27] = 32'b0000000_00111_00100_000_00000_0110011; // addi $t0, $0, 3 (error3)
  RegisterA[28] = 32'b0000000_01001_00010_000_00000_0110011; // addi $t1, $0, 3
  RegisterA[29] = 32'b0000000_01001_00000_000_00000_0110011;// 
  **/ 
end

assign InstructionOut = RegisterA[Address >> 2];

endmodule
